module demux_1to4_tb;
reg din;
reg [1:0] sel;
wire [3:0] dout;
demux_1to4 uut (.din(din), .sel(sel), .dout(dout));
initial begin
  $dumpfile("demux_1to4.vcd");
  $dumpvars(0, demux_1to4_tb);
  din = 1; sel = 2'b00;
  #10 sel = 2'b01;
  #10 sel = 2'b10;
  #10 sel = 2'b11;
  #10 $finish;
end
endmodule